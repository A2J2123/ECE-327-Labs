/***************************************************/
/* ECE 327: Digital Hardware Systems - Spring 2025 */
/* Lab 1 - Part 3                                  */
/* Testbench for ALU module                        */
/***************************************************/

`timescale 1ns/1ps

// Define the name of this testbench module. Since testbenches typically generate inputs and
// monitor outputs of the circuit being tested, they usually do not have any input/output ports.
module alu_tb ();

// Define any local parameters used in the testbench
localparam CLK_PERIOD = 8; // Clock period in nanoseconds
localparam DATAW = 4; // Bitwidth of ALU operands
localparam NUM_TESTS = 100; // Number of testcases generated by the testbench

// Declare logic signals for the circuit's inputs/outputs
logic clk_sig;
logic [DATAW-1:0] dataa_sig;
logic [DATAW-1:0] datab_sig;
logic [1:0] op_sig;
logic [2*DATAW-1:0] result_sig;

// Instantiate the design under test (dut), set the desired values of its parameters, and connect 
// its input/output ports to the declared signals.
alu # (
    .DATAW(DATAW)
) dut (
    .clk(clk_sig),
    .i_dataa(dataa_sig),
    .i_datab(datab_sig),
    .i_op(op_sig),
    .o_result(result_sig)
);

// Since the DUT tested here needs a clock signal, this initial block generates a clock signal with
// period 8ns and 50% duty cycle (i.e., 4ns high and 4ns low)
initial begin
    clk_sig = 1'b0;
    // The forever keyword means this keeps happening until the end of time (wait for half a clock
    // period, and flip its state)
    forever #(CLK_PERIOD/2) clk_sig = ~clk_sig; 
end

// The ALU circuit tested here has 3 inputs; 2x DATAW-bit inputs (operands) and 1x 2-bit input 
// (operation). It will be tedious to exhaustively test all possible input combinations, manually
// calculate their golden results, and visually verify the correctness of the produced outputs.
// Alternatively, we write code to randomly generate a number of test cases (NUM_TESTS), calculate
// the golden output using behavioral code, compare the produced outputs to these golden outputs,
// and automatically flag mismatches. Sometimes the golden outputs are even too complicated to be
// calculated in behavioral SystemVerilog. In such cases, we can implement a C++/Python software
// reference implementation which can generate test inputs and golden outputs and store them in a 
// file. Then, we can read these files in the SystemVerilog testbench to feed inputs to our DUT
// and verify its outputs.

// Declare variables used for test input and golden output generation
integer test_id; // Loop variable that goes from 0 to NUM_TESTS-1
integer correct_results; // Counter for correct outputs received from DUT
logic [2*DATAW-1:0] golden_result; // Golden result value to compare the output to

initial begin
    // Set time display format to be in 10^-9 sec, with 2 decimal places, and add " ns" suffix
    $timeformat(-9, 2, " ns");
    
    // Set all inputs to zeros and wait for 5 clock cycles
    dataa_sig = 'd0;
    datab_sig = 'd0;
    op_sig = 2'b00;
    correct_results = 0;
    #(5 * CLK_PERIOD);
    
    // Test the DUT using NUM_TESTS test cases
    for (test_id = 0; test_id < NUM_TESTS; test_id = test_id + 1) begin
        // For each test case, use Verilog system function $random to generate random inputs ...
        dataa_sig = $random;
        datab_sig = $random;
        op_sig = $random % 4; // Operation signal can be 0, 1, 2, or 3
        
        // ... and calculate the golden output for these inputs then wait 2 clock cycles
        if (op_sig == 2'b00) golden_result = 0;
        else if (op_sig == 2'b01) golden_result = dataa_sig << datab_sig;
        else if (op_sig == 2'b10) golden_result = signed'(dataa_sig) + signed'(datab_sig);
        else if (op_sig == 2'b11) golden_result = signed'(dataa_sig) - signed'(datab_sig);
        // We wait two clock cycles because we know the inputs and outputs are registered. Therefore,
        // the outputs of a set of inputs injected in cycle N will be produced in cycle N+2
        #(2*CLK_PERIOD);
        
        // Compare the DUT produced output to the golden output and display appropriate messages
        if (result_sig == golden_result) begin
            $write("[%0t] Correct Result! ", $time);
            correct_results = correct_results + 1;
        end else begin
            $write("[%0t] INCORRECT RESULT! ", $time);
        end
        case (op_sig)
            2'b00: $display("A=%b( %d)\t B=%b( %d)\t OP=RST\t\t Result=%b( %d)\t Golden=%b( %d)", dataa_sig, dataa_sig, datab_sig, datab_sig, result_sig, result_sig, golden_result, golden_result);
            2'b01: $display("A=%b( %d)\t B=%b( %d)\t OP=SHL\t\t Result=%b( %d)\t Golden=%b( %d)", dataa_sig, dataa_sig, datab_sig, datab_sig, result_sig, result_sig, golden_result, golden_result);
            2'b10: $display("A=%b(%d)\t B=%b(%d)\t OP=ADD\t\t Result=%b(%d)\t Golden=%b(%d)", signed'(dataa_sig), signed'(dataa_sig), signed'(datab_sig), signed'(datab_sig), signed'(result_sig), signed'(result_sig), signed'(golden_result), signed'(golden_result));
            2'b11: $display("A=%b(%d)\t B=%b(%d)\t OP=SUB\t\t Result=%b(%d)\t Golden=%b(%d)", signed'(dataa_sig), signed'(dataa_sig), signed'(datab_sig), signed'(datab_sig), signed'(result_sig), signed'(result_sig), signed'(golden_result), signed'(golden_result));
        endcase
    end
    
    // After all NUM_TESTS are completed, print the summary report and stop the simulation
    if (correct_results == NUM_TESTS) begin
        $display("Test PASSED! %d out of %d tests are matching golden outputs!", correct_results, NUM_TESTS);
    end else begin
        $display("Test FAILED! %d tests are not matching golden outputs!", NUM_TESTS - correct_results);
    end
    $stop;
end

endmodule